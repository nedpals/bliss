module main

import os